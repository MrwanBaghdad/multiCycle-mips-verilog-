module alu(in1,in2,aluop,out);
input [31:0]in1,in2;
output[31:0]out;
input []aluop;

case(aluop)

end module;