module mux3 (in1,in2,in3,chooser,out);

input [31:0] in1,in2,in3;
output [31:0] out;

